module ansi (
    input [7:0] a, d,
    output logic [7:0] q,
    input clk, reset_n
);

endmodule
