module Atop (a, b, c, d);

  localparam W = 16;

  input a;
  input [3:0] b, c;
  output [W-1:0] d;





endmodule
